`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    23:51:09 11/23/2014 
// Design Name: 
// Module Name:    camera_test_nexys2 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module camera_test_nexys2(
    input clk,
    input reset,
    input [7:0] JA,
    input [7:0] JB,
    input [7:0] JC,
    input [3:0] btn,
    output [7:0] Led,
    output [2:0] vgaRed,
    output [2:0] vgaGreen,
    output [1:0] vgaBlue,
    output Hsync,
    output Vsync,
    output clock_25mhz,
    inout sdiod,
    output sdioc,
    output xclk,
    output sccb_clk,
    output [6:0] seg,
    output dp,
    output [3:0] an
    );


endmodule

`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    23:51:09 11/23/2014 
// Design Name: 
// Module Name:    camera_test_nexys2 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module camera_test_nexys2(
    input clk,
    input reset,
    input [7:0] JA,
    input [7:0] JB,
    input [7:0] JC,
    input [3:0] btn,
    output [7:0] Led,
    output [2:0] vgaRed,
    output [2:0] vgaGreen,
    output [1:0] vgaBlue,
    output Hsync,
    output Vsync,
    output clock_25mhz,
    inout sdiod,
    output sdioc,
    output xclk,
    output sccb_clk,
    output [6:0] seg,
    output dp,
    output [3:0] an
    );


endmodule
