`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    09:38:46 12/08/2014 
// Design Name: 
// Module Name:    camera_sequencer 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module camera_sequencer(
	input clk,
	input start,
	output [31:0] beta_addr,
	output [31:0] beta_din,
	output [
    );


endmodule
