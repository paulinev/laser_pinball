library verilog;
use verilog.vl_types.all;
entity camera_read_tb is
end camera_read_tb;
