// top-level Verilog module for starter board (cjt, 10/05)
// * provides legit default values for all output pins (no floating tri-state!)
// * remember to comment out assignment to pins you will drive

module beta2demo(
     // clocks
     clock_50MHz, clock_socket,

     // 256k x 32 SRAM
     sram_a,sram_ce_b,sram_we_b,
     sram_io1,sram_ce1,sram_ub1,sram_lb1,
     sram_io2,sram_ce2,sram_ub2,sram_lb2,

     // I/O
     segment,an,sw,btn,led,
     vga_r,vga_g,vga_b,vga_hs,vga_vs,
     ps2_d,ps2_c,
     rs232_rxd,rs232_txd,rs232_rxd_a,rs232_txd_a,
     flash_d0,flash_oe,flash_rclk,

     // expansion connectors
     A1_4,A1_21,A1_22,
     A2_io,A2_db,A2_astb,A2_dstb,A2_write,A2_wait,A2_reset,
     B1_db,B1_adr,B1_we,B1_oe,B1_cs,B1_astb,B1_dstb,B1_write,B1_wait,B1_reset,B1_int
     );

   input clock_50MHz;
   input clock_socket;

   output [17:0] sram_a;
   output 	 sram_ce_b;
   output 	 sram_we_b;
   inout [15:0]  sram_io1;
   output 	 sram_ce1;
   output 	 sram_ub1;
   output 	 sram_lb1;
   inout [15:0]  sram_io2;
   output 	 sram_ce2;
   output 	 sram_ub2;
   output 	 sram_lb2;

   output [7:0]  segment;   // active low
   output [3:0]  an;        // active low
   input [7:0] 	 sw;
   input [3:0] 	 btn;
   output [7:0]  led;

   output 	 vga_r;
   output 	 vga_g;
   output 	 vga_b;
   output 	 vga_hs;
   output 	 vga_vs;

   inout 	 ps2_d;
   input 	 ps2_c;

   input 	 rs232_rxd;
   output 	 rs232_txd;
   input 	 rs232_rxd_a;
   output 	 rs232_txd_a;

   input 	 flash_d0;
   output 	 flash_oe;
   output 	 flash_rclk;

   inout 	 A1_4,A1_21,A1_22;

   inout [18:1]  A2_io;
   inout [7:0] 	 A2_db;
   inout 	 A2_astb;
   inout 	 A2_dstb;
   inout 	 A2_write;
   inout 	 A2_wait;
   inout 	 A2_reset;

   inout [7:0] 	 B1_db;
   inout [5:0] 	 B1_adr;
   inout 	 B1_we;
   inout 	 B1_oe;
   inout 	 B1_cs;
   inout 	 B1_astb;
   inout 	 B1_dstb;
   inout 	 B1_write;
   inout 	 B1_wait;
   inout 	 B1_reset;
   inout 	 B1_int;

   // SRAM pins
   assign sram_a = 18'h0;
   assign sram_ce_b = 1'b1;
   assign sram_we_b = 1'b1;
   assign sram_io1 = 18'h0;
   assign sram_ce1 = 1'b0;
   assign sram_ub1 = 1'b0;
   assign sram_lb1 = 1'b0;
   assign sram_io2 = 1'b0;
   assign sram_ce2 = 1'b0;
   assign sram_ub2 = 1'b0;
   assign sram_lb2 = 1'b0;

   // misc. I/O
   //assign segment = 8'hFF;   // active low
   //assign an = 4'hF;         // active low
   //assign led = 8'hAA;       // show it's us!!!
   //assign vga_r = 1'b0;
   //assign vga_g = 1'b0;
   //assign vga_b = 1'b0;
   //assign vga_hs = 1'b0;
   //assign vga_vs = 1'b0;
   assign ps2_d = 1'bz;
   assign rs232_txd = 1'b0;
   assign rs232_txd_a = 1'b0;
   assign flash_oe = 1'b1;
   assign flash_rclk = 1'b0;

   // expansion connectors
   assign A1_4 = 1'b0;
   assign A1_21 = 1'b0;
   assign A1_22 = 1'b0;
   assign A2_io = 18'h00000;
   assign A2_db = 8'h00;
   assign A2_astb = 1'b0;
   assign A2_dstb = 1'b0;
   assign A2_write = 1'b0;
   assign A2_wait = 1'b0;
   assign A2_reset = 1'b0;
   assign B1_db = 8'h00;
   assign B1_adr = 6'h00;
   assign B1_we = 1'b0;
   assign B1_oe = 1'b0;
   assign B1_cs = 1'b0;
   assign B1_astb = 1'b0;
   assign B1_dstb = 1'b0;
   assign B1_write = 1'b0;
   assign B1_wait = 1'b0;
   assign B1_reset = 1'b0;
   assign B1_int = 1'b0;

   //////////////////////////////////////////////////////////////////////
   //
   //  BETA2
   //
   //////////////////////////////////////////////////////////////////////

   wire clk,clk_300Hz;
   wire irq,irq_60Hz;
   wire [30:0] irq_addr;
  
   assign clk = clock_50MHz;

   wire power_on_reset;
   SRL16 reset_sr (.D(1'b0), .CLK(clk), .Q(power_on_reset),
		   .A0(1'b1), .A1(1'b1), .A2(1'b1), .A3(1'b1));
   defparam reset_sr.INIT = 16'hFFFF;

   wire user_reset;
   debounce dbreset(clk,btn[3],user_reset);

   wire reset = power_on_reset | user_reset;
   
   // make a Beta!
   wire mwe;
   reg [31:0] mdin;
   wire [31:0] ma,mdout,ramout,dpyout,ps2out;
   beta2 cpu(clk,reset,irq,irq_addr,ma,mdin,mdout,mwe);

   // decode memory address
   wire highmem = &ma[31:15];    // includes supervisor bit!
   wire sel_ram = !highmem;
   wire sel_dpy = highmem && ~ma[14];
   wire sel_60Hz = highmem && &ma[14:3] && ma[2];
   wire sel_ps2 = highmem && &ma[14:3] && ~ma[2];

   // remember what beta is trying to read
   reg [1:0] mdin_sel;
   reg rd_ps2;
   always @ (posedge clk) begin
      mdin_sel <= sel_dpy ? 2'd1 :
                  sel_ps2 ? 2'd2 :
                  2'd0;
      rd_ps2 <= !mwe && sel_ps2;
   end

   // select data to send back to beta
   always @ (mdin_sel or ramout or dpyout or ps2out)
     case (mdin_sel)
       default: mdin = ramout;
       2'd1: mdin = dpyout;
       2'd2: mdin = ps2out;
     endcase

   // program memory: up to 16K x 32
   // (memory module generated by betamem.py)
   lab9 mem(ma[15:2],clk,mdout,ramout,mwe & sel_ram);

   // 80x40 character display
   vga dpy(clk,vga_hs,vga_vs,{vga_r,vga_g,vga_b},irq_60Hz,sel_60Hz,
           mwe & sel_dpy,ma[11:2],mdout,dpyout);

   // ps2 interface
   ps2 kbd(clk,reset,clk_300Hz,ps2_c,ps2_d,
           rd_ps2,ps2out[7:0],ps2out[8],ps2out[9]);
   assign ps2out[31:10] = 0;

   // interrupts
   assign irq = ~ps2out[8] || irq_60Hz;
   assign irq_addr = ~ps2out[8] ? 12 : 8;
   assign led = {7'd0,irq};

   // show memory address in the 7-segments display
   segdisplay lights(clk,1'b1,ma[15:0],an,segment,clk_300Hz);

endmodule // beta2demo
