// 8x12 font memory for 128 chars
module xfont(addr,clk,row);
  input clk;
  input [10:0] addr;
  output [7:0] row;

  // font read-only memory: (128 * 12row/chars) x (8 bits/row)
  RAMB16_S9 font(.CLK(clk),.ADDR(addr),.DO(row),
                 .WE(1'b0),.EN(1'b1),.SSR(1'b0));
  defparam font.INIT_00 = 256'b00011000_00011000_00011000_00011000_00011000_00011000_00011000_00011000_11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam font.INIT_01 = 256'b00011000_00011000_00011000_00011000_00000000_00000000_00000000_00000000_00000000_11111000_11111000_00011000_00011000_00011000_00011000_00011000_00000000_00000000_00000000_00000000_00000000_11111111_11111111_00000000_00000000_00000000_00000000_00000000_00011000_00011000_00011000_00011000;
  defparam font.INIT_02 = 256'b00011000_00011000_00011000_00011000_00011000_11111000_11111000_00000000_00000000_00000000_00000000_00000000_00011000_00011000_00011000_00011000_00011000_00011111_00011111_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00011111_00011111_00011000;
  defparam font.INIT_03 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_11111111_10000001_10000001_10000001_10000001_10000001_10000001_10000001_10000001_10000001_10000001_11111111;
  defparam font.INIT_04 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam font.INIT_05 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam font.INIT_06 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam font.INIT_07 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam font.INIT_08 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam font.INIT_09 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam font.INIT_0A = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam font.INIT_0B = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam font.INIT_0C = 256'b00000000_00000000_00000000_00100100_01100110_01100110_01100110_00000000_00000000_00000000_00011000_00011000_00000000_00011000_00011000_00111100_00111100_00111100_00011000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam font.INIT_0D = 256'b01100010_00000000_00000000_00000000_00000000_00000000_00011000_00011000_01111100_00000110_00000110_00111100_01100000_01100000_00111110_00011000_00000000_00000000_00110110_00110110_01111111_00110110_00110110_00110110_01111111_00110110_00110110_00000000_00000000_00000000_00000000_00000000;
  defparam font.INIT_0E = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00110000_00011000_00011000_00011000_00000000_00000000_00000000_00111011_01101110_01100110_01111111_01111101_00111000_01101100_01101100_00111000_00000000_00000000_00000000_01000110_01100110_00110000_00011000_00001100_01100110;
  defparam font.INIT_0F = 256'b01100110_00111100_11111111_00111100_01100110_00000000_00000000_00000000_00000000_00000000_00110000_00011000_00001100_00000110_00000110_00000110_00001100_00011000_00110000_00000000_00000000_00000000_00000110_00001100_00011000_00110000_00110000_00110000_00011000_00001100_00000110_00000000;
  defparam font.INIT_10 = 256'b00000000_00000000_00000000_00000000_00000000_00110000_00011100_00011100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00011000_00011000_01111110_00011000_00011000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam font.INIT_11 = 256'b00000000_00000000_10000000_11000000_01100000_00110000_00011000_00001100_00000110_00000011_00000001_00000000_00000000_00000000_00011100_00011100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_01111110_00000000;
  defparam font.INIT_12 = 256'b00110000_00011000_00001100_00000110_01100011_01100011_00111110_00000000_00000000_00000000_01111110_00011000_00011000_00011000_00011000_00011000_01111000_00011000_00001000_00000000_00000000_00000000_00111110_01100011_01110011_01111011_01101011_01101111_01100111_01100011_00111110_00000000;
  defparam font.INIT_13 = 256'b01100000_01100000_01111110_00000000_00000000_00000000_00001111_00000110_00000110_01111111_01100110_00110110_00011110_00001110_00000110_00000000_00000000_00000000_00111110_01100011_00000011_00000011_00011110_00000011_00000011_01100011_00111110_00000000_00000000_00000000_01111111_01100011;
  defparam font.INIT_14 = 256'b00000000_00000000_00011000_00011000_00011000_00001100_00000110_00000011_00000011_01100011_01111111_00000000_00000000_00000000_00111100_01100110_01100110_01100110_01111100_01100000_01100000_00110000_00011100_00000000_00000000_00000000_00111100_01100110_00000110_00000110_00111100_01100000;
  defparam font.INIT_15 = 256'b00011100_00000000_00000000_00011100_00011100_00000000_00000000_00000000_00000000_00000000_00111000_00011000_00001100_00001100_00111110_01100110_01100110_01100110_00111100_00000000_00000000_00000000_00111100_01100110_01100110_01101110_00111100_00110110_01100110_01100110_00111100_00000000;
  defparam font.INIT_16 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000110_00001100_00011000_00110000_01100000_00110000_00011000_00001100_00000110_00000000_00000000_00011000_00001100_00011100_00011100_00000000_00000000_00011100_00011100_00000000_00000000_00000000_00000000_00000000_00000000_00011100;
  defparam font.INIT_17 = 256'b00000000_00000000_00001100_00001100_00000000_00001100_00001100_00000110_00000011_01100011_00111110_00000000_00000000_00000000_00110000_00011000_00001100_00000110_00000011_00000110_00001100_00011000_00110000_00000000_00000000_00000000_00000000_00000000_00000000_01111110_00000000_01111110;
  defparam font.INIT_18 = 256'b00110011_00110011_00111110_00110011_00110011_00110011_01111110_00000000_00000000_00000000_01100110_01100110_01100110_01111110_01100110_01100110_01100110_00111100_00011000_00000000_00000000_00000000_00111110_01100000_01100000_01101111_01101111_01101111_01100011_01100011_00111100_00000000;
  defparam font.INIT_19 = 256'b00110000_00110001_01111111_00000000_00000000_00000000_01111100_00110110_00110011_00110011_00110011_00110011_00110011_00110110_01111100_00000000_00000000_00000000_00011110_00110011_01100000_01100000_01100000_01100000_01100011_00110011_00011110_00000000_00000000_00000000_01111110_00110011;
  defparam font.INIT_1A = 256'b00000000_00000000_00011111_00110011_01100011_01100111_01100000_01100000_01100011_00110011_00011110_00000000_00000000_00000000_01111000_00110000_00110000_00110010_00111110_00110010_00110001_00110011_01111111_00000000_00000000_00000000_01111111_00110001_00110000_00110010_00111110_00110010;
  defparam font.INIT_1B = 256'b01100110_00000110_00000110_00000110_00000110_00000110_00001111_00000000_00000000_00000000_00111100_00011000_00011000_00011000_00011000_00011000_00011000_00011000_00111100_00000000_00000000_00000000_01100110_01100110_01100110_01100110_01111110_01100110_01100110_01100110_01100110_00000000;
  defparam font.INIT_1C = 256'b01111111_01110111_01100011_00000000_00000000_00000000_01111111_00110011_00110011_00110001_00110000_00110000_00110000_00110000_01111000_00000000_00000000_00000000_01110011_00110011_00110110_00110110_00111110_00110110_00110110_00110011_01110011_00000000_00000000_00000000_00111100_01100110;
  defparam font.INIT_1D = 256'b00000000_00000000_00011100_00110110_01100011_01100011_01100011_01100011_01100011_00110110_00011100_00000000_00000000_00000000_01100011_01100011_01100111_01101111_01111111_01111011_01110011_01100011_01100011_00000000_00000000_00000000_01100011_01100011_01100011_01100011_01100011_01101011;
  defparam font.INIT_1E = 256'b00110011_00110110_00111110_00110011_00110011_00110011_01111110_00000000_00000000_00000000_00001111_00000110_00111110_01101111_01100111_01100011_01100011_00110110_00011100_00000000_00000000_00000000_01111000_00110000_00110000_00110000_00111110_00110011_00110011_00110011_01111110_00000000;
  defparam font.INIT_1F = 256'b01100110_01100110_01100110_00000000_00000000_00000000_00111100_00011000_00011000_00011000_00011000_00011000_00011000_01011010_01111110_00000000_00000000_00000000_00111100_01100110_01100110_00001100_00111000_01100000_01100110_01100110_00111100_00000000_00000000_00000000_01110011_00110011;
  defparam font.INIT_20 = 256'b00000000_00000000_00110110_00110110_01101011_01101011_01100011_01100011_01100011_01100011_01100011_00000000_00000000_00000000_00011000_00111100_01100110_01100110_01100110_01100110_01100110_01100110_01100110_00000000_00000000_00000000_00111100_01100110_01100110_01100110_01100110_01100110;
  defparam font.INIT_21 = 256'b00110001_00110000_00011000_00001100_00001100_01100111_01111111_00000000_00000000_00000000_00111100_00011000_00011000_00011000_00111100_01100110_01100110_01100110_01100110_00000000_00000000_00000000_01100110_01100110_01100110_00111100_00011000_00111100_01100110_01100110_01100110_00000000;
  defparam font.INIT_22 = 256'b00000110_00000110_00011110_00000000_00000000_00000000_00000001_00000011_00000110_00001100_00011000_00110000_01100000_01000000_00000000_00000000_00000000_00000000_00011110_00011000_00011000_00011000_00011000_00011000_00011000_00011000_00011110_00000000_00000000_00000000_01111111_01100011;
  defparam font.INIT_23 = 256'b00000000_01111111_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_01100011_00110110_00011100_00001000_00000000_00000000_00011110_00000110_00000110_00000110_00000110_00000110;
  defparam font.INIT_24 = 256'b00110011_00110011_00111110_00110000_00110000_00110000_01110000_00000000_00000000_00000000_00111011_01100110_01100110_00111110_00000110_00111100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00110000_01100000_01100000;
  defparam font.INIT_25 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00111011_01100110_01100110_01100110_01100110_00111110_00000110_00000110_00001110_00000000_00000000_00000000_00111100_01100110_01100000_01100000_01100110_00111100_00000000_00000000_00000000_00000000_00000000_00000000_01101110_00110011;
  defparam font.INIT_26 = 256'b00111100_01100110_00000110_00111110_01100110_01100110_01100110_00111011_00000000_00000000_00000000_00000000_00000000_00000000_00111100_00011000_00011000_00011000_00111110_00011000_00011000_00011011_00001110_00000000_00000000_00000000_00111100_01100110_01100000_01111110_01100110_00111100;
  defparam font.INIT_27 = 256'b00000110_00000110_00000110_00011110_00000000_00000110_00000110_00000000_00000000_00000000_00111111_00001100_00001100_00001100_00001100_00111100_00000000_00001100_00001100_00000000_00000000_00000000_01110011_00110011_00110011_00110011_00111011_00110110_00110000_00110000_01100000_00000000;
  defparam font.INIT_28 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00111111_00001100_00001100_00001100_00001100_00001100_00001100_00001100_00111100_00000000_00000000_00000000_01110011_00110011_00110110_00111100_00110110_00110011_00110000_00110000_01110000_00000000_00111100_01100100_01100110_00000110;
  defparam font.INIT_29 = 256'b00000000_00000000_00111100_01100110_01100110_01100110_01100110_00111100_00000000_00000000_00000000_00000000_00000000_00000000_01100110_01100110_01100110_01100110_01100110_01111100_00000000_00000000_00000000_00000000_00000000_00000000_01100011_01101011_01101011_01101011_01101011_01111110;
  defparam font.INIT_2A = 256'b00110000_00111011_00110111_01110110_00000000_00000000_00000000_00000000_00001111_00000110_00111110_01100110_01100110_01100110_01100110_00111011_00000000_00000000_00000000_00000000_01111000_00110000_00111110_00110011_00110011_00110011_00110011_01101110_00000000_00000000_00000000_00000000;
  defparam font.INIT_2B = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00011100_00110110_00110000_00110000_00110000_01111110_00110000_00010000_00000000_00000000_00000000_00000000_00111100_01100110_00001100_00110000_01100110_00111100_00000000_00000000_00000000_00000000_00000000_00000000_01111000_00110000;
  defparam font.INIT_2C = 256'b00000000_00000000_00110110_00110110_01101011_01101011_01100011_01100011_00000000_00000000_00000000_00000000_00000000_00000000_00011000_00111100_01100110_01100110_01100110_01100110_00000000_00000000_00000000_00000000_00000000_00000000_00111011_01100110_01100110_01100110_01100110_01100110;
  defparam font.INIT_2D = 256'b00011000_00000110_01000011_01111111_00000000_00000000_00000000_00000000_01111000_00001100_00000110_00011110_00110011_00110011_00110011_00110011_00000000_00000000_00000000_00000000_00000000_00000000_01100011_00110110_00011100_00011100_00110110_01100011_00000000_00000000_00000000_00000000;
  defparam font.INIT_2E = 256'b00011000_00011000_01110000_00000000_00000000_00000000_00011000_00011000_00011000_00011000_00000000_00011000_00011000_00011000_00011000_00000000_00000000_00000000_00000111_00001100_00001100_00011000_00110000_00011000_00001100_00001100_00000111_00000000_00000000_00000000_01111111_01100001;
  defparam font.INIT_2F = 256'b00000000_00000000_01111110_01111110_01111110_01111110_01111110_01111110_01111110_01111110_01111110_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_11001110_11011010_01110011_00000000_00000000_00000000_01110000_00011000_00011000_00001100_00000110_00001100;
  defparam font.INIT_30 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam font.INIT_31 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam font.INIT_32 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam font.INIT_33 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam font.INIT_34 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam font.INIT_35 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam font.INIT_36 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam font.INIT_37 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam font.INIT_38 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam font.INIT_39 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam font.INIT_3A = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam font.INIT_3B = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam font.INIT_3C = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam font.INIT_3D = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam font.INIT_3E = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam font.INIT_3F = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;

endmodule