library verilog;
use verilog.vl_types.all;
entity camera_save_with_read_tb is
end camera_save_with_read_tb;
