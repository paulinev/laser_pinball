`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    21:22:45 12/02/2014 
// Design Name: 
// Module Name:    my_ic2 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module my_ic2(
	input wire clk,
	input wire [7:0] din,
	input wire start,
	input wire stop,
	input wire sda_i,
	output wire sda_o,
	output wire sda_o_en,
	
	
	inout wire scl
    );
	 
	 


endmodule
