// single-port read/write memory initialized with lab9 code
module lab9(addr,clk,din,dout,we);
  input [13:0] addr;     // up to 16K locations
  input clk;             // memory has internal address regs
  input [31:0] din;      // appears after rising clock edge
  output [31:0] dout;    // written at rising clock edge
  input we;              // enables write port

  // we're using 1833 out of 2048 locations
  RAMB16_S9 m0(.CLK(clk),.ADDR(addr[10:0]),.DI(din[7:0]),.DO(dout[7:0]),.WE(we),.EN(1'b1),.SSR(1'b0),.DIP(1'b0));
  defparam m0.INIT_00 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00100001_00000011_00000100_00101100_00110101;
  defparam m0.INIT_01 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_10011000_00000000_00000000_00000000_00000000_00000000;
  defparam m0.INIT_02 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m0.INIT_03 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m0.INIT_04 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m0.INIT_05 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m0.INIT_06 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m0.INIT_07 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m0.INIT_08 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m0.INIT_09 = 256'b01011000_01010100_01010000_01001100_01001000_01000100_01000000_00111100_00111000_00110100_00110000_00101100_00101000_00100100_00100000_00011100_00011000_00010100_11111111_00101110_01110010_01101110_01100101_01110000_01010101_10001000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m0.INIT_0A = 256'b11001100_11001100_11001100_11001100_11001100_11001100_11001100_11001100_11001100_11001100_11001100_10110000_11001100_00000000_01001100_00000010_00011010_11111100_10010100_10001100_10001000_10000100_10000000_01111100_01111000_01110100_01110000_01101100_01101000_01100100_01100000_01011100;
  defparam m0.INIT_0B = 256'b01110100_01101100_00100000_00110010_00011000_11111100_00000000_01101001_01110010_01101001_01100111_01001001_00111011_11001100_11001100_11001100_11001100_11001100_11001100_11001100_11001100_11001100_11001100_11001100_11001100_11001100_11001100_11001100_11001100_11001100_11001100_11001100;
  defparam m0.INIT_0C = 256'b01110100_01110000_01101100_01101000_01100100_01100000_01011100_01011000_01010100_01010000_01001100_01001000_01000100_01000000_00111100_00111000_00110100_00110000_00101100_00101000_00100100_00100000_00011100_00011000_00010100_11111111_00101110_00100001_00101011_00010001_11111100_00100000;
  defparam m0.INIT_0D = 256'b11000111_11100100_00010100_11100100_11101011_11100100_00000000_11010000_01000000_00101100_01001100_11101000_00110000_00111100_00101000_00000000_11000100_00000010_00000111_11111100_11011011_00001001_10001100_00000100_10001100_00000000_10001100_10001000_10000100_10000000_01111100_01111000;
  defparam m0.INIT_0E = 256'b00011101_00010101_00001101_01100110_01010101_01001110_01000101_01000110_00111110_00111101_00110110_00101110_00100101_00100110_00011110_00010110_00001110_00000111_01111000_00001001_00000001_00001010_10000011_00001011_00000011_00001100_00000100_00000110_00000101_01110110_00000000_00000000;
  defparam m0.INIT_0F = 256'b01001001_01000001_00111010_00110001_00110010_00101010_00100001_00100010_00011010_01011010_01010010_01001100_01001011_01000010_00111011_00110011_00110100_00101011_00100011_00011011_00011100_01011101_01011011_01010100_01001101_01000100_01000011_00111100_00110101_00101100_00101101_00100100;
  defparam m0.INIT_10 = 256'b00010100_00100000_01011001_00100000_00010010_00000000_00000000_11110010_00000000_00000010_11110000_11110110_11100000_11111111_00000000_00011100_00011000_00010100_00000100_00000000_11111000_00011100_00011000_00010100_00000100_00000000_01110010_01101011_01110100_01110101_00101001_01001010;
  defparam m0.INIT_11 = 256'b00000000_00000101_00000000_00000111_00000000_00000000_00000100_11010010_11010011_11100100_00000000_11111111_00001000_00000001_00000000_00000100_00001000_00000000_11111001_00000100_00000010_00000000_11100001_11111111_00000000_00001000_11100101_00010011_01011000_00100000_00010001_00100000;
  defparam m0.INIT_12 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00110001_00111111_00010100_00110100_10001100_01100110_10001100_00111000_00000111_00010100_11111011_00000000_11111111_11000010_00000100_00000000_00000011_00000100_00000000_00000001_00000000_00000011;
  defparam m0.INIT_13 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_01011000_01111000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m0.INIT_14 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_01101000_10001000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m0.INIT_15 = 256'b00010100_11001100_01011000_00000001_11001100_01111100_11001100_00001101_11001100_00010100_11111100_00000100_01011000_10001000_10011100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m0.INIT_16 = 256'b00110000_00110000_00101100_00101100_00101000_00101000_00100100_00100100_00100000_00100000_00011100_00011100_00011000_00011000_00010100_00010100_00010000_00010000_00001100_00001100_00001000_00001000_00000100_00000100_00000000_00000000_00000000_11111100_11111100_00011000_00010100_00000101;
  defparam m0.INIT_17 = 256'b01110000_01110000_01101100_01101100_01101000_01101000_01100100_01100100_01100000_01100000_01011100_01011100_01011000_01011000_01010100_01010100_01010000_01010000_01001100_01001100_01001000_01001000_01000100_01000100_01000000_01000000_00111100_00111100_00111000_00111000_00110100_00110100;
  defparam m0.INIT_18 = 256'b01001000_01000100_01000000_00111100_00111000_00110100_00110000_00101100_00101000_00100100_00100000_00011100_00011000_00010100_00010100_00000000_00010100_00000010_00000000_00011000_00000001_00011000_00010100_11111100_00000100_00000000_00000010_00000000_01111000_01111000_01110100_01110100;
  defparam m0.INIT_19 = 256'b01010000_00110000_11111100_10000000_00000100_00000000_00000000_00000100_00000000_10010100_01010001_01111111_01010011_10000001_10010100_10001100_10001000_10000100_10000000_01111100_01111000_01110100_01110000_01101100_01101000_01100100_01100000_01011100_01011000_01010100_01010000_01001100;
  defparam m0.INIT_1A = 256'b00001101_10000000_01010000_00000011_00001010_11111100_00000100_11111100_00000100_11111100_00000100_00110000_00110011_00000000_00000001_00000000_00110111_00000000_00000001_01011010_00000000_01011100_00100001_01101000_01001000_00000000_01011000_01111000_00000100_00100000_00000000_00011100;
  defparam m0.INIT_1B = 256'b11111100_11111100_11111100_01010000_11111100_11111100_00000001_00000000_00000000_00000000_11111111_00000000_00000000_00000000_00000011_00000011_11111111_11111100_00000100_00001111_00001010_00110000_11111100_10000000_00000100_00000000_11111011_00110000_00000100_00000000_01010000_00000000;
  defparam m0.INIT_1C = 256'b00000100_00011100_00000000_00001000_11111100_00000100_11111100_00000100_11111100_00000100_11111100_00000100_01000110_01000101_01000100_01000011_01000010_01000001_00111001_00111000_00110111_00110110_00110101_00110100_00110011_00110010_00110001_00110000_00000000_11111100_11111100_11111100;
  defparam m0.INIT_1D = 256'b00000000_11111100_00000100_11111100_00000100_11111100_00000100_11111100_00000100_00000000_11111100_11111100_00000000_00000100_00000000_11111100_00000100_00000000_11111100_11111100_11111100_11111100_11111100_11111100_11111100_11111100_11111000_00000001_10110001_00010000_00000010_00001111;
  defparam m0.INIT_1E = 256'b11110100_11111100_00000100_00001010_01101110_00101100_01110000_01110100_01010011_00000001_00000001_01010100_00000000_11111100_11111100_11111100_11111100_11111100_11111100_11111100_11111100_00000000_11110110_11111010_00000001_00001000_10001111_00000101_01111111_00000100_00000100_00000000;
  defparam m0.INIT_1F = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_11111010_00000100_11100110_00001010_01101011_00000000_01110100_11111000_00001010_00000100_00000000_11110000_00000010_11111111_00000011_01110100_00111110_00000001_00000100_10011100_00001010_00000001_11111100_11111100_00000101;
  defparam m0.INIT_20 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m0.INIT_21 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m0.INIT_22 = 256'b00000000_00000000_11100100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m0.INIT_23 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m0.INIT_24 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m0.INIT_25 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m0.INIT_26 = 256'b11111100_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m0.INIT_27 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_01011001_00000011_01010101_00000101_01001111_00000111_01001001_00001001_01000101_00001011_01000001_00000000_11111100_11111100_00100000_00000001_01100001_00000011_01111010;
  defparam m0.INIT_28 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m0.INIT_29 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m0.INIT_2A = 256'b01100100_01111100_00000000_01110100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m0.INIT_2B = 256'b00000100_11111100_00000100_00000000_11111100_11111100_11111100_11111100_11111100_11111100_00000110_11100111_11111100_00000100_01101000_00000000_00000001_01100100_00000001_11011000_00000010_01101000_11111100_11111100_00000101_11110111_11111100_00000100_11111100_00000100_11111100_00000100;
  defparam m0.INIT_2C = 256'b00100000_00000101_01001010_11100000_00000000_10000100_00000000_11111100_11111100_11111100_11111100_11111100_11111100_00000110_11001100_11111100_00000100_01101100_00000000_00000001_01100100_00000001_11011000_00000010_01101100_11111100_11111100_00000101_11011000_11111100_00000100_11111100;
  defparam m0.INIT_2D = 256'b00000000_00000000_00000000_11011110_11111100_11111100_00000110_00011011_11111100_00000100_11100101_00001010_00000010_00000000_01000001_00000001_11111010_00000010_00000100_00000000_00000100_00000000_00000000_00000000_11111100_00100000_11010111_00000010_11111000_00000100_00000000_00000111;
  defparam m0.INIT_2E = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m0.INIT_2F = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m0.INIT_30 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m0.INIT_31 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_11110100_00000000;
  defparam m0.INIT_32 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m0.INIT_33 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m0.INIT_34 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m0.INIT_35 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_11111011_00000111_10011100_00000001_10011100_00000000_00000000;
  defparam m0.INIT_36 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m0.INIT_37 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m0.INIT_38 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m0.INIT_39 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m0.INIT_3A = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m0.INIT_3B = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m0.INIT_3C = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m0.INIT_3D = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m0.INIT_3E = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m0.INIT_3F = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  RAMB16_S9 m1(.CLK(clk),.ADDR(addr[10:0]),.DI(din[15:8]),.DO(dout[15:8]),.WE(we),.EN(1'b1),.SSR(1'b0),.DIP(1'b0));
  defparam m1.INIT_00 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000011_00000001_00000011;
  defparam m1.INIT_01 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m1.INIT_02 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m1.INIT_03 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m1.INIT_04 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m1.INIT_05 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m1.INIT_06 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m1.INIT_07 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m1.INIT_08 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m1.INIT_09 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_11111111_00101110_01110101_01110100_01100100_01100101_01101110_00000010_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m1.INIT_0A = 256'b00000101_00000101_00000101_00000101_00000101_00000101_00000101_00000101_00000101_00000101_00000101_00000110_00000101_00000000_00000101_00000000_00000000_11111111_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m1.INIT_0B = 256'b01101001_01101111_01100001_00000010_00000010_11111111_00000000_01101111_01110101_01101110_01100001_01101100_00000010_00000101_00000101_00000101_00000101_00000101_00000101_00000101_00000101_00000101_00000101_00000101_00000101_00000101_00000101_00000101_00000101_00000101_00000101_00000101;
  defparam m1.INIT_0C = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_11111111_00101110_00100000_00000010_00000010_11111111_00110000;
  defparam m1.INIT_0D = 256'b11111111_00000110_00000000_00000110_11111111_00000110_00000000_00001100_00001101_00001101_00001001_00000110_00001001_00001001_00001101_00000000_00000110_00000000_00000000_11111111_11111111_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m1.INIT_0E = 256'b01110111_01110001_00001001_00001000_00111101_00101101_00110000_00111001_00111000_00110111_00110110_00110101_00110100_00110011_00110010_00110001_01100000_10001100_10001011_10001010_10001001_10001000_10000111_10000110_10000101_10000100_10000011_10000010_10000001_00110011_00000000_00000000;
  defparam m1.INIT_0F = 256'b00101110_00101100_01101101_01101110_01100010_01110110_01100011_01111000_01111010_00001010_00100111_00111011_01101100_01101011_01101010_01101000_01100111_01100110_01100100_01110011_01100001_01011100_01011101_01011011_01110000_01101111_01101001_01110101_01111001_01110100_01110010_01100101;
  defparam m1.INIT_10 = 256'b00000000_00000000_00000000_00000000_00000000_00000111_00000111_11111111_00000111_00000000_00000000_11111111_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_11111111_00000000_00000000_00000000_00000000_00000000_10010011_10010010_10010001_10010000_00100000_00101111;
  defparam m1.INIT_11 = 256'b00000010_00000000_00000001_00000000_00000100_00000100_00000111_11111111_11111111_00000110_00010000_00000000_00000000_00000000_00000111_00000111_00000000_00000000_11111111_00000000_00000000_00010000_11111111_00000000_00000000_00000111_11111111_00000000_00000000_00000000_00000000_00000000;
  defparam m1.INIT_12 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_11111111_00000001_00000000_11111111_00000000_00000001_00000000_11111111_00000001_00000000_11111111_00000000_11111111_11111111_00000111_00000000_00000000_00000111_00010000_00000000_00001000_00000000;
  defparam m1.INIT_13 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00001111_00010001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m1.INIT_14 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00010110_00011000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m1.INIT_15 = 256'b00000000_00001010_00001001_00000000_00001010_00000000_00001010_00000000_00001010_00000000_11111111_00000000_00001001_00011010_00011010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m1.INIT_16 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_11111111_11111111_00001100_00001100_00000000;
  defparam m1.INIT_17 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m1.INIT_18 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00001100_00000000_00001100_00000000_11111111_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m1.INIT_19 = 256'b00001101_10001100_11111111_10001100_00000000_00000000_10000000_00000111_00000111_00000000_11111110_11111111_11111110_11111111_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m1.INIT_1A = 256'b00000000_10001100_00001101_00000000_00000000_11111111_00000000_11111111_00000000_11111111_00000000_10001100_11111110_00000000_00000000_00000000_11111110_00000000_00000000_11111110_00000000_11111110_00000000_01100101_01101001_00000000_00001111_00010001_00000000_00001101_00000000_00001101;
  defparam m1.INIT_1B = 256'b11111111_11111111_11111111_00001101_11111111_11111111_00000000_00000000_00010000_00010000_11111111_00000000_00010000_00010000_00000000_00000000_00000000_11111111_00000000_00000000_00000000_10001100_11111111_10001100_00000000_00000000_11111111_10001100_00000000_00000000_00000000_10000000;
  defparam m1.INIT_1C = 256'b00000000_00000000_11111000_00000000_11111111_00000000_11111111_00000000_11111111_00000000_11111111_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_11111111_11111111_11111111;
  defparam m1.INIT_1D = 256'b11111000_11111111_00000000_11111111_00000000_11111111_00000000_11111111_00000000_00000000_11111111_11111111_11111000_00000000_11111000_11111111_00000000_00000000_11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111_00000000_11111111_00001110_00000000_00000000;
  defparam m1.INIT_1E = 256'b11111111_11111111_00000000_00001010_01101011_00100000_01101001_00100000_01110100_00000000_00000000_00001111_00000000_11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111000_11111111_11111111_00000000_00000000_11111111_00000000_00000000_00000000_00000000_00000000;
  defparam m1.INIT_1F = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_11111111_00000000_11111111_00000000_00000001_00000000_00010001_11111111_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00010001_00100000_00000000_00000000_00011100_00000000_00000000_11111111_11111111_00000000;
  defparam m1.INIT_20 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m1.INIT_21 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m1.INIT_22 = 256'b00000000_00000000_00001111_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m1.INIT_23 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m1.INIT_24 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m1.INIT_25 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m1.INIT_26 = 256'b11111111_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m1.INIT_27 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_11111111_11111111_00000000_00000000_00000000_00000000_00000000;
  defparam m1.INIT_28 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m1.INIT_29 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m1.INIT_2A = 256'b00000000_00010101_00000000_00010101_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m1.INIT_2B = 256'b00000000_11111111_00000000_00000000_11111111_11111111_11111111_11111111_11111111_11111111_00000000_11111111_11111111_00000000_00010101_00000000_00000000_00000000_00000000_00010011_00000000_00010101_11111111_11111111_00000000_11111111_11111111_00000000_11111111_00000000_11111111_00000000;
  defparam m1.INIT_2C = 256'b00000000_00000000_11111111_11111111_11111000_00011000_00000000_11111111_11111111_11111111_11111111_11111111_11111111_00000000_11111111_11111111_00000000_00010101_00000000_00000000_00000000_00000000_00010011_00000000_00010101_11111111_11111111_00000000_11111111_11111111_00000000_11111111;
  defparam m1.INIT_2D = 256'b00000000_00000000_00000000_11111111_11111111_11111111_00000000_11111110_11111111_00000000_11111111_00000000_00000000_11111000_01011001_00000000_11111111_00000000_00000000_00000000_00000000_00101000_11111000_11111000_11111111_00000000_11111111_00000000_11111111_00000000_00000000_00000000;
  defparam m1.INIT_2E = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m1.INIT_2F = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m1.INIT_30 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m1.INIT_31 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00010110_00000000;
  defparam m1.INIT_32 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m1.INIT_33 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m1.INIT_34 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m1.INIT_35 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_11111111_00000000_00011100_00000000_00011100_00000000_00000000;
  defparam m1.INIT_36 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m1.INIT_37 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m1.INIT_38 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m1.INIT_39 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m1.INIT_3A = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m1.INIT_3B = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m1.INIT_3C = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m1.INIT_3D = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m1.INIT_3E = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m1.INIT_3F = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  RAMB16_S9 m2(.CLK(clk),.ADDR(addr[10:0]),.DI(din[23:16]),.DO(dout[23:16]),.WE(we),.EN(1'b1),.SSR(1'b0),.DIP(1'b0));
  defparam m2.INIT_00 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_11111111_11111111_11111111_11111111_11111111;
  defparam m2.INIT_01 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m2.INIT_02 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m2.INIT_03 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m2.INIT_04 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m2.INIT_05 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m2.INIT_06 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m2.INIT_07 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m2.INIT_08 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m2.INIT_09 = 256'b00111111_00011111_11111111_11011111_10111111_10011111_01111111_01011111_00111111_00011111_11111111_11011111_10111111_10011111_01111111_01011111_00111111_00011111_11111111_00101110_01110000_01100101_00100000_01100011_01100101_10011111_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m2.INIT_0A = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_11100000_00000000_00000000_00000000_00011110_10111111_11011111_10111111_10011111_01111111_01011111_00111111_00011111_11111111_11011111_10111111_10011111_01111111_01011111;
  defparam m2.INIT_0B = 256'b01101111_01100011_01110100_10011111_10011111_00011110_00000000_01101110_01100011_01110011_01101100_01101100_10011111_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m2.INIT_0C = 256'b00011111_11111111_11011111_10111111_10011111_01111111_01011111_00111111_00011111_11111111_11011111_10111111_10011111_01111111_01011111_00111111_00011111_11111111_11011111_10111111_10011111_01111111_01011111_00111111_00011111_11111111_00101110_00101110_10011111_10011111_00011110_01111000;
  defparam m2.INIT_0D = 256'b11111111_11111111_00011111_00011111_11100000_00011111_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_11100000_00000000_00000000_00000000_00011110_11111111_10011111_00011111_00000000_00011111_11111110_11011111_10111111_10011111_01111111_01011111_00111111;
  defparam m2.INIT_0E = 256'b01010111_01010001_00001001_00001000_00101011_01011111_00101001_00101000_00101010_00100110_01011110_00100101_00100100_00100011_01000000_00100001_01111110_10001100_10001011_10001010_10001001_10001000_10000111_10000110_10000101_10000100_10000011_10000010_10000001_00110011_00000000_00000000;
  defparam m2.INIT_0F = 256'b00111110_00111100_01001101_01001110_01000010_01010110_01000011_01011000_01011010_00001010_00100010_00111010_01001100_01001011_01001010_01001000_01000111_01000110_01000100_01010011_01000001_01111100_01111101_01111011_01010000_01001111_01001001_01010101_01011001_01010100_01010010_01000101;
  defparam m2.INIT_10 = 256'b00100000_11100001_00100000_11100001_00100000_11111111_01011111_11111111_00011111_11100001_00100000_11100001_00100000_00000000_11111110_01011111_00111111_00011111_11100001_00100000_00011111_01011111_00111111_00011111_11011110_00000000_10010011_10010010_10010001_10010000_00100000_00111111;
  defparam m2.INIT_11 = 256'b00011111_11111111_00011111_11111111_00011111_01000010_01011111_11100010_11111111_00111111_00100001_00100001_00100001_11100000_00000010_01011111_00100001_00100001_11111111_00100001_11100010_01000000_11100010_01000010_01000001_00111111_11100010_11100001_00100000_11100001_00100000_11100001;
  defparam m2.INIT_12 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_11111111_10011111_00011111_11111111_00011111_10011111_00011111_11111111_10011111_00011111_11111111_00100001_00000000_11111111_00111111_00100001_11100010_00111111_00011111_11111111_00011111_11111111;
  defparam m2.INIT_13 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m2.INIT_14 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m2.INIT_15 = 256'b00111111_00011111_00011111_11100001_00100000_00000000_00011111_10011111_00111111_00011111_10011101_10111101_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m2.INIT_16 = 256'b01000001_01000000_01000001_01000000_01000001_01000000_01000001_01000000_01000001_01000000_01000001_01000000_01000001_01000000_01000001_01000000_01000001_01000000_01000001_01000000_01000001_01000000_01000001_01000000_01000001_01000000_11111100_10111101_10011101_00011111_00011111_10011111;
  defparam m2.INIT_17 = 256'b01000001_01000000_01000001_01000000_01000001_01000000_01000001_01000000_01000001_01000000_01000001_01000000_01000001_01000000_01000001_01000000_01000001_01000000_01000001_01000000_01000001_01000000_01000001_01000000_01000001_01000000_01000001_01000000_01000001_01000000_01000001_01000000;
  defparam m2.INIT_18 = 256'b10111111_10011111_01111111_01011111_00111111_00011111_11111111_11011111_10111111_10011111_01111111_01011111_00111111_00011111_00011111_11111110_00011111_11100000_00000000_00011111_00000000_00011111_00011111_11111111_11011110_00000000_00000000_11111100_01000001_01000000_01000001_01000000;
  defparam m2.INIT_19 = 256'b00011111_00011111_11100001_00100000_00000000_11100000_00011111_11111111_11111111_10111111_11111111_10011111_11111111_10011111_10111111_11011111_10111111_10011111_01111111_01011111_00111111_00011111_11111111_11011111_10111111_10011111_01111111_01011111_00111111_00011111_11111111_11011111;
  defparam m2.INIT_1A = 256'b11100010_01000001_00111111_11100010_01000000_01011101_10111101_00111101_10111101_00011101_10111101_11111111_11111111_00000011_00000000_00000011_11111111_00000011_00000000_11100000_00000011_11111111_00000000_01110010_00100000_11111110_11011111_10111111_00100000_00111111_00100000_00111111;
  defparam m2.INIT_1B = 256'b00111101_10111101_01011101_00111111_10111101_01111101_00100001_01000001_01000000_01000011_01100011_01000001_01100011_00000000_01000010_01000001_01111111_01111101_10111101_11100010_01000000_00111111_11100010_01000001_00100001_11100001_11100010_01000001_00100001_01000001_01000001_00111111;
  defparam m2.INIT_1C = 256'b00100001_00000001_00100000_01011111_01011101_10111101_00111101_10111101_00011101_10111101_10011101_10111101_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_11111100_10111101_00011101_10111101;
  defparam m2.INIT_1D = 256'b00100000_01111101_10111101_01011101_10111101_00111101_10111101_10011101_10111101_11111100_10111101_00011101_10000000_10011111_00011100_00011101_10111101_11111100_10111101_10011101_10111101_00011101_10111101_00111101_10111101_01011101_11100010_01000010_10011111_00000000_00000000_00000000;
  defparam m2.INIT_1E = 256'b01100000_01111101_10111101_00000000_01111001_01000010_01101110_01110100_01100001_00000000_00000000_00000000_11111100_10111101_10011101_10111101_00111101_10111101_01011101_10111101_01111101_00000001_11111111_11100011_01100011_01000010_10011111_11100000_00000010_01111111_00100001_01000001;
  defparam m2.INIT_1F = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_11111111_01000010_11100001_00100000_10011111_00000010_01011111_11100001_00100000_01100011_00000011_10011111_00000000_00000000_00000000_01111111_00000000_00000000_00000000_00011111_00000000_00000000_10111101_01111101_00000000;
  defparam m2.INIT_20 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m2.INIT_21 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m2.INIT_22 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m2.INIT_23 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m2.INIT_24 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m2.INIT_25 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m2.INIT_26 = 256'b00111101_10111101_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m2.INIT_27 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_11111100_00111111_11100001_00100000_11100001_00100000_11100001_00100000_11100001_00100000_11100001_00100000_11100001_00100000_11111100_10111101_00111101_00000000_11100001_00100000_11100001_00100000;
  defparam m2.INIT_28 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m2.INIT_29 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m2.INIT_2A = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m2.INIT_2B = 256'b10111101_00111101_10111101_11111100_10111101_00111101_10111101_01011101_10111101_01111101_00000000_01100000_01111101_10111101_00111111_00111111_11100010_01000001_00100001_00000010_01000001_00111111_10111101_01111101_00000000_01100000_01111101_10111101_01011101_10111101_00111101_10111101;
  defparam m2.INIT_2C = 256'b00100000_11100001_10011111_10011111_10101001_00111111_11111100_10111101_00111101_10111101_01011101_10111101_01111101_00000000_01100000_01111101_10111101_00111111_00111111_11100010_01000001_00100001_00000010_01000001_00111111_10111101_01111101_00000000_01100000_01111101_10111101_01011101;
  defparam m2.INIT_2D = 256'b00000000_00000000_00000000_11111111_10111101_01111101_00000000_01100000_01111101_10111101_11100000_00000011_00000000_00000011_00000000_00000000_11111111_00000000_10000100_00000100_11100001_00100100_10001001_01100000_11100001_00100000_10011111_00000000_11111111_10100101_00000101_11100001;
  defparam m2.INIT_2E = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m2.INIT_2F = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m2.INIT_30 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m2.INIT_31 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m2.INIT_32 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m2.INIT_33 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m2.INIT_34 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m2.INIT_35 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_11111111_00000000_00011111_00000000_00011111_00000000_00000000;
  defparam m2.INIT_36 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m2.INIT_37 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m2.INIT_38 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m2.INIT_39 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m2.INIT_3A = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m2.INIT_3B = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m2.INIT_3C = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m2.INIT_3D = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m2.INIT_3E = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m2.INIT_3F = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  RAMB16_S9 m3(.CLK(clk),.ADDR(addr[10:0]),.DI(din[31:24]),.DO(dout[31:24]),.WE(we),.EN(1'b1),.SSR(1'b0),.DIP(1'b0));
  defparam m3.INIT_00 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_01110111_01110111_01110111_01110111_01110111;
  defparam m3.INIT_01 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m3.INIT_02 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m3.INIT_03 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m3.INIT_04 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m3.INIT_05 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m3.INIT_06 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m3.INIT_07 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m3.INIT_08 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m3.INIT_09 = 256'b01100110_01100110_01100101_01100101_01100101_01100101_01100101_01100101_01100101_01100101_01100100_01100100_01100100_01100100_01100100_01100100_01100100_01100100_01110111_00000000_01110100_01110010_01101001_01110100_01111000_01110111_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m3.INIT_0A = 256'b10000000_10000000_10000000_10000000_10000000_10000000_10000000_10000000_10000000_10000000_10000000_10000000_10000000_01101111_01100000_11110000_11110100_01100000_01100011_01100111_01100111_01100111_01100111_01100111_01100111_01100111_01100110_01100110_01100110_01100110_01100110_01100110;
  defparam m3.INIT_0B = 256'b01101110_01100001_00100000_01110111_01110111_01100000_00000000_00100000_01110100_01110100_00100000_01100101_01110111_10000000_10000000_10000000_10000000_10000000_10000000_10000000_10000000_10000000_10000000_10000000_10000000_10000000_10000000_10000000_10000000_10000000_10000000_10000000;
  defparam m3.INIT_0C = 256'b01100011_01100010_01100010_01100010_01100010_01100010_01100010_01100010_01100010_01100001_01100001_01100001_01100001_01100001_01100001_01100001_01100001_01100000_01100000_01100000_01100000_01100000_01100000_01100000_01100000_01110111_00000000_00101110_01110111_01110111_11000100_00000000;
  defparam m3.INIT_0D = 256'b01110111_01100111_01100100_01100000_01110111_01100000_00000000_10000000_10000000_10000000_10000000_10000000_10000000_10000000_10000000_01101111_01100000_11110000_11100000_01100000_01110111_01110111_01100100_11000100_01100000_01101111_01100011_01100011_01100011_01100011_01100011_01100011;
  defparam m3.INIT_0E = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m3.INIT_0F = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m3.INIT_10 = 256'b11010000_01111011_11010000_01111011_11010000_01100111_01100000_01110111_01100100_01110111_11010000_01111011_11010000_11100000_01101111_01100000_01100000_01100000_01110111_11100000_01100000_01100100_01100100_01100100_11000111_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m3.INIT_11 = 256'b11000000_01110111_11000000_01110111_11000000_11100000_01100000_01110111_01110111_01100100_10100100_11100000_11110100_01110111_11100000_01100000_11110100_01100000_01110111_11000000_01111011_10010000_01110111_11100000_01100000_11000000_01111011_01111011_11010000_01111011_11010000_01111011;
  defparam m3.INIT_12 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_01110111_01110111_01100000_01110111_01100100_01110111_01100000_01110111_01110111_01100000_01110111_10100000_11101000_01110111_01100100_10100100_01111011_01100000_11000000_01110111_11000000_01110111;
  defparam m3.INIT_13 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m3.INIT_14 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m3.INIT_15 = 256'b11000000_01100100_11000000_01111011_11010100_11000000_01100000_01110111_01100000_11000000_01100111_11000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m3.INIT_16 = 256'b01100100_01100000_01100100_01100000_01100100_01100000_01100100_01100000_01100100_01100000_01100100_01100000_01100100_01100000_01100100_01100000_01100100_01100000_01100100_01100000_01100100_01100000_01100100_01100000_01100100_01100000_01101111_11000011_01100011_01100100_01100000_01110111;
  defparam m3.INIT_17 = 256'b01100100_01100000_01100100_01100000_01100100_01100000_01100100_01100000_01100100_01100000_01100100_01100000_01100100_01100000_01100100_01100000_01100100_01100000_01100100_01100000_01100100_01100000_01100100_01100000_01100100_01100000_01100100_01100000_01100100_01100000_01100100_01100000;
  defparam m3.INIT_18 = 256'b01100101_01100101_01100101_01100101_01100101_01100101_01100100_01100100_01100100_01100100_01100100_01100100_01100100_01100100_01100000_01101111_01100000_01111011_11010100_01100100_11000100_01100000_01100100_01100011_11000111_00000000_00000000_01101111_01100100_01100000_01100100_01100000;
  defparam m3.INIT_19 = 256'b01100100_11000000_01111011_11010100_11000000_01100111_11000000_01100111_01100111_01100011_01110111_01110111_01110111_01110111_01100011_01100111_01100111_01100111_01100111_01100111_01100111_01100111_01100110_01100110_01100110_01100110_01100110_01100110_01100110_01100110_01100101_01100101;
  defparam m3.INIT_1A = 256'b01111011_11010100_01100000_01111011_11010000_01100100_11000011_01100100_11000011_01100100_11000011_11111111_01110111_01100100_11000000_01100000_01110111_01100100_11000100_01110111_01100000_01110111_00000000_01100101_01110100_01101111_11000011_11000011_01100100_01100000_01100100_01100000;
  defparam m3.INIT_1B = 256'b01100000_11000011_01100000_01100100_11000011_01100000_11000000_01100100_10100100_10100000_11101000_01100000_10110000_10110000_11110000_11100000_11000000_01100100_11000011_01111011_11010000_11000000_01111011_11010100_11000000_01100111_01111011_11010100_11000000_01100100_01100000_11000000;
  defparam m3.INIT_1C = 256'b11110000_11111000_10000000_11000000_01100100_11000011_01100100_11000011_01100100_11000011_01100111_11000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_01101111_11000011_01100000_11000011;
  defparam m3.INIT_1D = 256'b10000000_01100100_11000011_01100100_11000011_01100100_11000011_01100111_11000011_01101111_11000011_01100000_10000011_01110111_10000000_01100100_11000011_01101111_11000011_01100011_11000011_01100000_11000011_01100000_11000011_01100000_01111011_11000100_01110111_01100000_11110000_11100000;
  defparam m3.INIT_1E = 256'b01111100_01100100_11000011_00000000_00101110_01110101_01100111_01111001_01110010_00000100_00000000_00000000_01101111_11000011_01100011_11000011_01100000_11000011_01100000_11000011_01100000_10000000_01110111_01111011_11000100_11111000_01110111_01110111_11100000_11000000_11000000_01100000;
  defparam m3.INIT_1F = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_01110111_11000000_01111011_11010000_01110111_01100000_01100000_01110111_11010000_11000000_01100100_01110111_00000100_11100000_00000100_01100000_00000000_00000100_00000100_01100000_00000000_00000100_11000011_01100000_00000100;
  defparam m3.INIT_20 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m3.INIT_21 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m3.INIT_22 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m3.INIT_23 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m3.INIT_24 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m3.INIT_25 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m3.INIT_26 = 256'b01100100_11000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m3.INIT_27 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_01101111_11000000_01111011_11010000_01111011_11010000_01111011_11010000_01111011_11010000_01111011_11010000_01111011_11010000_01101111_11000011_01100000_11000100_01111011_11010100_01110111_11011000;
  defparam m3.INIT_28 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m3.INIT_29 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m3.INIT_2A = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m3.INIT_2B = 256'b11000011_01100100_11000011_01101111_11000011_01100000_11000011_01100000_11000011_01100000_00000100_01111100_01100100_11000011_01100100_11000000_01110111_11010000_11000000_01100100_11110000_01100000_11000011_01100000_00000100_01111100_01100100_11000011_01100100_11000011_01100100_11000011;
  defparam m3.INIT_2C = 256'b11011000_01111011_01110111_01110111_10000000_01100001_01101111_11000011_01100000_11000011_01100000_11000011_01100000_00000100_01111100_01100100_11000011_01100100_11000000_01110111_11010000_11000000_01100000_11110000_01100000_11000011_01100000_00000100_01111100_01100100_11000011_01100100;
  defparam m3.INIT_2D = 256'b00000000_00000000_00000000_01110111_11000011_01100000_00000100_01111100_01100100_11000011_01110111_11010000_00000100_10000000_00000000_00000100_01110111_00000100_11000000_01100000_01111011_10010000_10000000_10000000_01110111_11011000_01110111_00000100_01110111_11000000_01100100_01111011;
  defparam m3.INIT_2E = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m3.INIT_2F = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m3.INIT_30 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m3.INIT_31 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m3.INIT_32 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m3.INIT_33 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m3.INIT_34 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m3.INIT_35 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_01110111_00000100_01100100_11000000_01100000_00000000_00000000;
  defparam m3.INIT_36 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m3.INIT_37 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m3.INIT_38 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m3.INIT_39 = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m3.INIT_3A = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m3.INIT_3B = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m3.INIT_3C = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m3.INIT_3D = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m3.INIT_3E = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
  defparam m3.INIT_3F = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;

endmodule